`ifndef RKV_WATCHDOG_SEQ_LIB_SVH
`define RKV_WATCHDOG_SEQ_LIB_SVH

`include "rkv_watchdog_element_sequences.svh" //why comp element before base_virtual 
`include "rkv_watchdog_base_virtual_sequence.sv"

`include "rkv_watchdog_integration_virt_seq.sv"
`include "rkv_watchdog_apbacc_virt_seq.sv"
`include "rkv_watchdog_regacc_virt_seq.sv"
`include "rkv_watchdog_countdown_virt_seq.sv"
`include "rkv_watchdog_resen_virt_seq.sv"
`include "rkv_watchdog_disable_intr_virt_seq.sv"
`include "rkv_watchdog_lock_virt_seq.sv"
`include "rkv_watchdog_reload_virt_seq.sv"

`endif 
