`ifndef RKV_WATCHDOG_TESTS_SVH
`define RKV_WATCHDOG_TESTS_SVH

`include "rkv_watchdog_base_test.sv"
`include "rkv_watchdog_integration_test.sv"
`include "rkv_watchdog_apbacc_test.sv"
`include "rkv_watchdog_regacc_test.sv"
`include "rkv_watchdog_countdown_test.sv"
`include "rkv_watchdog_resen_test.sv"
`include "rkv_watchdog_disable_intr_test.sv"
`include "rkv_watchdog_lock_test.sv"
`include "rkv_watchdog_reload_test.sv"

`endif // RKV_WATCHDOG_TESTS_SVH
