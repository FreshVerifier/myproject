`ifndef RKV_WATCHDOG_COV_SVH
`define RKV_WATCHDOG_COV_SVH

`include "rkv_watchdog_cov.sv"

`endif //RKV_WATCHDOG_COV_SV
